DUT (.clk_in(intf.clk_in),
.free_l2clk(intf.free_l2clk	),
.active_clk(intf.active_clk	),
.rst_l(intf.rst_l	),
.dec_i0_decode_d(intf.dec_i0_decode_d	),
.exu_flush_final(intf.exu_flush_final	),
.dec_tlu_i0_commit_cmt(intf.dec_tlu_i0_commit_cmt	),
.dec_tlu_flush_err_wb(intf.dec_tlu_flush_err_wb	),
.dec_tlu_flush_noredir_wb(intf.dec_tlu_flush_noredir_wb	),
.exu_flush_path_final(intf.exu_flush_path_final	),
.dec_tlu_mrac_ff(intf.dec_tlu_mrac_ff	),
.dec_tlu_fence_i_wb(intf.dec_tlu_fence_i_wb	),
.dec_tlu_flush_leak_one_wb(intf.dec_tlu_flush_leak_one_wb	),
.dec_tlu_bpred_disable(intf.dec_tlu_bpred_disable	),
.dec_tlu_core_ecc_disable(intf.dec_tlu_core_ecc_disable	),
.dec_tlu_force_halt(intf.dec_tlu_force_halt	),
.ifu_axi_awvalid(intf.ifu_axi_awvalid	),
.ifu_axi_awid(intf.ifu_axi_awid	),
.ifu_axi_awaddr(intf.ifu_axi_awaddr	),
.ifu_axi_awregion(intf.ifu_axi_awregion	),
.ifu_axi_awlen(intf.ifu_axi_awlen	),
.ifu_axi_awsize(intf.ifu_axi_awsize	),
.ifu_axi_awburst(intf.ifu_axi_awburst	),
.ifu_axi_awlock(intf.ifu_axi_awlock	),
.ifu_axi_awcache(intf.ifu_axi_awcache	),
.ifu_axi_awprot(intf.ifu_axi_awprot	),
.ifu_axi_awqos(intf.ifu_axi_awqos	),
.ifu_axi_wvalid(intf.ifu_axi_wvalid	),
.ifu_axi_wdata(intf.ifu_axi_wdata	),
.ifu_axi_wstrb(intf.ifu_axi_wstrb	),
.ifu_axi_wlast(intf.ifu_axi_wlast	),
.ifu_axi_bready(intf.ifu_axi_bready	),
.ifu_axi_arvalid(intf.ifu_axi_arvalid	),
.ifu_axi_arready(intf.ifu_axi_arready	),
.ifu_axi_arid(intf.ifu_axi_arid	),
.ifu_axi_araddr(intf.ifu_axi_araddr	),
.ifu_axi_arregion(intf.ifu_axi_arregion	),
.ifu_axi_arlen(intf.ifu_axi_arlen	),
.ifu_axi_arsize(intf.ifu_axi_arsize	),
.ifu_axi_arburst(intf.ifu_axi_arburst	),
.ifu_axi_arlock(intf.ifu_axi_arlock	),
.ifu_axi_arcache(intf.ifu_axi_arcache	),
.ifu_axi_arprot(intf.ifu_axi_arprot	),
.ifu_axi_arqos(intf.ifu_axi_arqos	),
.ifu_axi_rvalid(intf.ifu_axi_rvalid	),
.ifu_axi_rready(intf.ifu_axi_rready	),
.fu_axi_rid(intf.fu_axi_rid	),
.ifu_axi_rdata(intf.ifu_axi_rdata	),
.ifu_axi_rresp(intf.ifu_axi_rresp	),
.ifu_bus_clk_en(intf.ifu_bus_clk_en	),
.dma_iccm_req(intf.dma_iccm_req	),
.dma_mem_addr(intf.dma_mem_addr	),
.dma_mem_sz(intf.dma_mem_sz	),
.dma_mem_write(intf.dma_mem_write	),
.dma_mem_wdata(intf.dma_mem_wdata	),
.dma_mem_tag(intf.dma_mem_tag	),
.dma_iccm_stall_any(intf.dma_iccm_stall_any	),
.iccm_dma_ecc_error(intf.iccm_dma_ecc_error	),
.iccm_dma_rvalid(intf.iccm_dma_rvalid	),
.iccm_dma_rdata(intf.iccm_dma_rdata	),
.iccm_dma_rtag(intf.iccm_dma_rtag	),
.iccm_ready(intf.iccm_ready	),
.ifu_pmu_instr_aligned(intf.ifu_pmu_instr_aligned	),
.ifu_pmu_fetch_stall(intf.ifu_pmu_fetch_stall	),
.ifu_ic_error_start(intf.ifu_ic_error_start	),
.ic_rw_addr(intf.ic_rw_addr	),
.ic_wr_en(intf.ic_wr_en	),
.ic_rd_en(intf.ic_rd_en	),
.ic_wr_data(intf.ic_wr_data	),
.ic_rd_data(intf.ic_rd_data	),
.ic_debug_rd_data(intf.ic_debug_rd_data	),
.ictag_debug_rd_data(intf.ictag_debug_rd_data	),
.ic_debug_wr_data(intf.ic_debug_wr_data	),
.ifu_ic_debug_rd_data(intf.ifu_ic_debug_rd_data	),
.ic_eccerr(intf.ic_eccerr	),
.ic_parerr(intf.ic_parerr	),
.ic_premux_data(intf.ic_premux_data	),
.ic_sel_premux_data(intf.ic_sel_premux_data	),
.ic_debug_addr(intf.ic_debug_addr	),
.ic_debug_rd_en(intf.ic_debug_rd_en	),
.ic_debug_wr_en(intf.ic_debug_wr_en	),
.ic_debug_tag_array(intf.ic_debug_tag_array	),
.ic_debug_way(intf.ic_debug_way	),
.ic_tag_valid(intf.ic_tag_valid	),
.ic_rd_hit(intf.ic_rd_hit	),
.ic_tag_perr(intf.ic_tag_perr	),
.iccm_rw_addr(intf.iccm_rw_addr	),
.iccm_wren(intf.iccm_wren	),
.iccm_rden(intf.iccm_rden	),
.iccm_wr_data(intf.iccm_wr_data	),
.iccm_wr_size(intf.iccm_wr_size	),
.iccm_rd_data(intf.iccm_rd_data	),
.iccm_rd_data_ecc(intf.iccm_rd_data_ecc	),
.ifu_iccm_rd_ecc_single_err(intf.ifu_iccm_rd_ecc_single_err	),
.ifu_pmu_ic_miss(intf.ifu_pmu_ic_miss	),
.ifu_pmu_ic_hit(intf.ifu_pmu_ic_hit	),
.ifu_pmu_bus_error(intf.ifu_pmu_bus_error	),
.ifu_pmu_bus_busy(intf.ifu_pmu_bus_busy	),
.ifu_pmu_bus_trxn(intf.ifu_pmu_bus_trxn	),
.ifu_i0_icaf(intf.ifu_i0_icaf	),
.ifu_i0_icaf_type(intf.ifu_i0_icaf_type	),
.ifu_i0_valid(intf.ifu_i0_valid	),
.ifu_i0_icaf_second(intf.ifu_i0_icaf_second	),
.ifu_i0_dbecc(intf.ifu_i0_dbecc	),
.iccm_dma_sb_error(intf.iccm_dma_sb_error	),
.ifu_i0_instr(intf.ifu_i0_instr	),
.ifu_i0_pc(intf.ifu_i0_pc	),
.ifu_i0_pc4(intf.ifu_i0_pc4	),
.ifu_miss_state_idle(intf.ifu_miss_state_idle	),
.i0_brp(intf.i0_brp	),
.ifu_i0_bp_index(intf.ifu_i0_bp_index	),
.ifu_i0_bp_fghr(intf.ifu_i0_bp_fghr	),
.ifu_i0_bp_btag(intf.ifu_i0_bp_btag	),
.ifu_i0_fa_index(intf.ifu_i0_fa_index	),
.exu_mp_pkt(intf.exu_mp_pkt	),
.exu_mp_eghr(intf.exu_mp_eghr	),
.exu_mp_fghr(intf.exu_mp_fghr	),
.exu_mp_index(intf.exu_mp_index	),
.exu_mp_btag(intf.exu_mp_btag	),
.dec_tlu_br0_r_pkt(intf.dec_tlu_br0_r_pkt	),
.exu_i0_br_fghr_r(intf.exu_i0_br_fghr_r	),
.exu_i0_br_index_r(intf.exu_i0_br_index_r	),
.dec_fa_error_index(intf.dec_fa_error_index	),
.dec_tlu_flush_lower_wb(intf.dec_tlu_flush_lower_wb	),
.ifu_i0_cinst(intf.ifu_i0_cinst	),
.dec_tlu_ic_diag_pkt(intf.dec_tlu_ic_diag_pkt	),
.ifu_ic_debug_rd_data_valid(intf.ifu_ic_debug_rd_data_valid	),
.iccm_buf_correct_ecc(intf.iccm_buf_correct_ecc	),
.iccm_correction_state(intf.iccm_correction_state	),
.scan_mode(intf.scan_mode	);